`ifndef __ALU_SV
`define __ALU_SV

module alu
    import common::*;
    import pipes::*;(
        
    );

    /* TODO: implement your ALU here. */

endmodule

`endif
