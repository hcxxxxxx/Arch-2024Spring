`ifndef __FORWARD_SV
`define __FORWARD_SV

module forward
    import common::*;
    import pipes::*;(
        input logic clk, reset
    );

    //useless

endmodule

`endif
