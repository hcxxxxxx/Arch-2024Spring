`ifndef __HAZARD_SV
`define __HAZARD_SV

module hazard
    import common::*;
    import pipes::*;(
        
    );

    

endmodule

`endif
